module top();
  initial 
    begin
      $display("hello world!");
    end
endmodule
